module comp5(input x,input y,input z,output w); 

 assign w = (x & z)|(x & y);
 
endmodule

 
